module sevenseg
(
	input [3:0] in,
	output [11:0] out //The data sheets are 1 indexed
);

case(in)
	0: out = 12'b011001001011;
	1: out = 12'b000001001000;
	2: out = 12'b010001010011;
	3: out = 12'b010001011010;
	4: out = 12'b001001011000;
	5: out = 12'b011000011010;
	6: out = 12'b011000011111;
	7: out = 12'b011001001000;
	8: out = 12'b011001011011;
	9: out = 12'b011001011010;
	3'hA: out = 12'b011001011001;
	3'hB: out = 12'b001000011011;
	3'hC: out = 12'b011000000011;
	3'hD: out = 12'b000001011011;
	3'hE: out = 12'b011000010011;
	3'hF: out = 12'b011000010001;
endcase
endmodule

/*

Digit 	gfedcba 	abcdefg 	a(11) 	b(7) 	c(4) 	d(2) 	e(1) 	f(10) 	g(5)
0 	0×3F 	0×7E 				1 		1 		1 		1 		1 		1 		0
1 	0×06 	0×30 				0 		1 		1 		0 		0 		0 		0
2 	0×5B 	0×6D 				1 		1 		0 		1 		1 		0 		1
3 	0×4F 	0×79 				1 		1 		1 		1 		0 		0 		1
4 	0×66 	0×33 				0 		1 		1 		0 		0 		1 		1
5 	0×6D 	0×5B 				1 		0 		1 		1 		0 		1 		1
6 	0×7D 	0×5F 				1 		0 		1 		1 		1 		1 		1
7 	0×07 	0×70 				1 		1 		1 		0 		0 		1 		0
8 	0×7F 	0×7F 				1 		1 		1 		1 		1 		1 		1
9 	0×6F 	0×7B 				1 		1 		1 		1 		0 		1 		1
A 	0×77 	0×77 				1 		1 		1 		0 		1 		1 		1
b 	0×7C 	0×1F 				0 		0 		1 		1 		1 		1 		1
C 	0×39 	0×4E 				1 		0 		0 		1 		1 		1 		0
d 	0×5E 	0×3D 				0 		1 		1 		1 		1 		0 		1
E 	0×79 	0×4F 				1 		0 		0 		1 		1 		1 		1
F 	0×71 	0×47 				1 		0 		0 		0 		1 		1 		1

*/
