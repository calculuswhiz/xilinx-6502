module dev_zero (
    input   [7:0] datain,
    output  [7:0] dataout
);

dataout = 8'h00;

endmodule
